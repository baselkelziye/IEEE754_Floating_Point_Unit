module clz(
    input  [23:0] in,   // 24-bit input
    output [4:0] count  // 5-bit output (since max leading zeros = 24)
);

    reg [4:0] cnt;

    always @(*) begin
        casez (in)
            24'b1??????????????????????? : cnt = 5'd0;
            24'b01?????????????????????? : cnt = 5'd1;
            24'b001????????????????????? : cnt = 5'd2;
            24'b0001???????????????????? : cnt = 5'd3;
            24'b00001??????????????????? : cnt = 5'd4;
            24'b000001?????????????????? : cnt = 5'd5;
            24'b0000001????????????????? : cnt = 5'd6;
            24'b00000001???????????????? : cnt = 5'd7;
            24'b000000001??????????????? : cnt = 5'd8;
            24'b0000000001?????????????? : cnt = 5'd9;
            24'b00000000001????????????? : cnt = 5'd10;
            24'b000000000001???????????? : cnt = 5'd11;
            24'b0000000000001??????????? : cnt = 5'd12;
            24'b00000000000001?????????? : cnt = 5'd13;
            24'b000000000000001????????? : cnt = 5'd14;
            24'b0000000000000001???????? : cnt = 5'd15;
            24'b00000000000000001??????? : cnt = 5'd16;
            24'b000000000000000001?????? : cnt = 5'd17;
            24'b0000000000000000001????? : cnt = 5'd18;
            24'b00000000000000000001???? : cnt = 5'd19;
            24'b000000000000000000001??? : cnt = 5'd20;
            24'b0000000000000000000001?? : cnt = 5'd21;
            24'b00000000000000000000001? : cnt = 5'd22;
            24'b000000000000000000000001 : cnt = 5'd23;
            default                      : cnt = 5'd24; // All zeros
        endcase
    end

    assign count = cnt;

endmodule
